library ieee;
use ieee.std_logic_1164.all;

entity random_gen is
  port (
    Clock : in std_logic 
  );
end random_gen;

architecture rtl of random_gen is
begin

end rtl;