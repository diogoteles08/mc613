library ieee;
use ieee.std_logic_1164.all;

entity type_proc is
  port (
    Clock : in std_logic
  );
end type_proc;

architecture rtl of type_proc is
begin

end rtl;