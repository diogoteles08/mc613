library ieee;
use ieee.std_logic_1164.all;

entity screen_proc is
  port (
    Clock : in std_logic;
 
  );
end screen_proc;

architecture rtl of screen_proc is
begin

end rtl;