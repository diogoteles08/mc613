library ieee;
use ieee.std_logic_1164.all;

entity word_gen is
  port (
    Clock : in std_logic;
 
  );
end word_gen;

architecture rtl of word_gen is

begin

end rtl;