library ieee;
use ieee.std_logic_1164.all;

entity clock_parser is
  port (
    Clock : in std_logic 
  );
end clock_parser;

architecture rtl of clock_parser is
begin

end rtl;