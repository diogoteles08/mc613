-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition"
-- CREATED		"Thu May 17 20:31:26 2018"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY CPU IS 
	PORT
	(
		clock :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		IO_IN :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		Pc_Ld :  OUT  STD_LOGIC;
		IR_Ld :  OUT  STD_LOGIC;
		Pc_Inc :  OUT  STD_LOGIC;
		ALU_2_DBus :  OUT  STD_LOGIC;
		DM_Rd :  OUT  STD_LOGIC;
		DM_Wr :  OUT  STD_LOGIC;
		PC_Ld_En :  OUT  STD_LOGIC;
		Reg_2_IO :  OUT  STD_LOGIC;
		IO_2_Reg :  OUT  STD_LOGIC;
		Reg_Wr :  OUT  STD_LOGIC;
		Stat_Wr :  OUT  STD_LOGIC;
		DM_2_DBus :  OUT  STD_LOGIC;
		DBus :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		IM_address :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		IM_instruction_out :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		instruction :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		IO_OUT :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		RSource1 :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		RSource2 :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		stat_CVNZ :  OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END CPU;

ARCHITECTURE bdf_type OF CPU IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT mux_0
	PORT(data : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 result : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF mux_0: COMPONENT IS true;
ATTRIBUTE noopt OF mux_0: COMPONENT IS true;

COMPONENT alu
GENERIC (WORDSIZE : INTEGER
			);
	PORT(A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Op : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 Z : OUT STD_LOGIC;
		 C : OUT STD_LOGIC;
		 V : OUT STD_LOGIC;
		 N : OUT STD_LOGIC;
		 F : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT memory
GENERIC (BITS_OF_ADDR : INTEGER;
			MIF_FILE : STRING;
			WORDSIZE : INTEGER
			);
	PORT(clock : IN STD_LOGIC;
		 we : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 datain : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 dataout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pc
GENERIC (increment : INTEGER;
			WORDSIZE : INTEGER
			);
	PORT(clock : IN STD_LOGIC;
		 clear : IN STD_LOGIC;
		 PC_Ld : IN STD_LOGIC;
		 PC_Inc : IN STD_LOGIC;
		 DATA_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT bank
GENERIC (WORDSIZE : INTEGER
			);
	PORT(WR_EN : IN STD_LOGIC;
		 RD_EN : IN STD_LOGIC;
		 clear : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 DATA_IN : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 RD_ADDR1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 RD_ADDR2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 WR_ADDR : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 DATA_OUT1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 DATA_OUT2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT reg
GENERIC (WORDSIZE : INTEGER
			);
	PORT(clock : IN STD_LOGIC;
		 load : IN STD_LOGIC;
		 clear : IN STD_LOGIC;
		 datain : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 dataout : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT uc
	PORT(clear : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 instruction : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 IR_Ld : OUT STD_LOGIC;
		 PC_Inc : OUT STD_LOGIC;
		 ALU_2_DBus : OUT STD_LOGIC;
		 DM_Rd : OUT STD_LOGIC;
		 DM_Wr : OUT STD_LOGIC;
		 PC_Ld_En : OUT STD_LOGIC;
		 Reg_2_IO : OUT STD_LOGIC;
		 IO_2_Reg : OUT STD_LOGIC;
		 Reg_Wr : OUT STD_LOGIC;
		 Stat_Wr : OUT STD_LOGIC;
		 DM_2_DBus : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	addr :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	ALU_2_DBus_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	C :  STD_LOGIC;
SIGNAL	DM_2_DBus_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	DM_Rd_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	DM_Wr_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	gdfx_temp0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	gnd :  STD_LOGIC;
SIGNAL	instruction_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	IO_2_Reg_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	IR_Ld_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	N :  STD_LOGIC;
SIGNAL	Pc_Inc_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	Pc_Ld_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	PC_Ld_En_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	preir :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	Reg_2_IO_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	Reg_Wr_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	Rs1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	Rs2 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	stat :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	Stat_Wr_ALTERA_SYNTHESIZED :  STD_LOGIC;
SIGNAL	V :  STD_LOGIC;
SIGNAL	vcc :  STD_LOGIC;
SIGNAL	Z :  STD_LOGIC;
SIGNAL	zeros :  STD_LOGIC_VECTOR(27 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;

SIGNAL	GDFX_TEMP_SIGNAL_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	GDFX_TEMP_SIGNAL_0 :  STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN 

GDFX_TEMP_SIGNAL_1 <= (zeros(27 DOWNTO 0) & C & V & N & Z);
GDFX_TEMP_SIGNAL_0 <= (zeros(5 DOWNTO 0) & instruction_ALTERA_SYNTHESIZED(25 DOWNTO 0));


b2v_ALU : alu
GENERIC MAP(WORDSIZE => 32
			)
PORT MAP(A => Rs1,
		 B => Rs2,
		 Op => instruction_ALTERA_SYNTHESIZED(27 DOWNTO 26),
		 Z => Z,
		 C => C,
		 V => V,
		 N => N,
		 F => SYNTHESIZED_WIRE_4);


b2v_D_Memory : memory
GENERIC MAP(BITS_OF_ADDR => 10,
			MIF_FILE => "dmemory.mif",
			WORDSIZE => 32
			)
PORT MAP(clock => clock,
		 we => DM_Wr_ALTERA_SYNTHESIZED,
		 address => Rs1(9 DOWNTO 0),
		 datain => Rs2,
		 dataout => SYNTHESIZED_WIRE_5);


b2v_I_Memory : memory
GENERIC MAP(BITS_OF_ADDR => 10,
			MIF_FILE => "fibonacci.mif",
			WORDSIZE => 32
			)
PORT MAP(clock => clock,
		 we => gnd,
		 address => addr(9 DOWNTO 0),
		 dataout => preir);




SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_0 XOR instruction_ALTERA_SYNTHESIZED(28);


b2v_inst13 : pc
GENERIC MAP(increment => 1,
			WORDSIZE => 32
			)
PORT MAP(clock => clock,
		 clear => reset,
		 PC_Ld => Pc_Ld_ALTERA_SYNTHESIZED,
		 PC_Inc => Pc_Inc_ALTERA_SYNTHESIZED,
		 DATA_IN => GDFX_TEMP_SIGNAL_0,
		 DATA_OUT => addr);


b2v_inst4 : bank
GENERIC MAP(WORDSIZE => 32
			)
PORT MAP(WR_EN => Reg_Wr_ALTERA_SYNTHESIZED,
		 RD_EN => vcc,
		 clear => reset,
		 clock => clock,
		 DATA_IN => gdfx_temp0,
		 RD_ADDR1 => instruction_ALTERA_SYNTHESIZED(20 DOWNTO 16),
		 RD_ADDR2 => instruction_ALTERA_SYNTHESIZED(15 DOWNTO 11),
		 WR_ADDR => instruction_ALTERA_SYNTHESIZED(25 DOWNTO 21),
		 DATA_OUT1 => Rs1,
		 DATA_OUT2 => Rs2);


SYNTHESIZED_WIRE_6 <= DM_Rd_ALTERA_SYNTHESIZED OR DM_2_DBus_ALTERA_SYNTHESIZED;


SYNTHESIZED_WIRE_2 <= instruction_ALTERA_SYNTHESIZED(28) AND instruction_ALTERA_SYNTHESIZED(27) AND instruction_ALTERA_SYNTHESIZED(26);


SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2;


Pc_Ld_ALTERA_SYNTHESIZED <= PC_Ld_En_ALTERA_SYNTHESIZED AND SYNTHESIZED_WIRE_3;


b2v_IR : reg
GENERIC MAP(WORDSIZE => 32
			)
PORT MAP(clock => clock,
		 load => IR_Ld_ALTERA_SYNTHESIZED,
		 clear => reset,
		 datain => preir,
		 dataout => instruction_ALTERA_SYNTHESIZED);


b2v_mux4to1 : mux_0
PORT MAP(data => stat(3 DOWNTO 0),
		 sel => instruction_ALTERA_SYNTHESIZED(27 DOWNTO 26),
		 result => SYNTHESIZED_WIRE_0);

zeros <= (gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd);



b2v_Status : reg
GENERIC MAP(WORDSIZE => 32
			)
PORT MAP(clock => clock,
		 load => Stat_Wr_ALTERA_SYNTHESIZED,
		 clear => reset,
		 datain => GDFX_TEMP_SIGNAL_1,
		 dataout => stat);


PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(31) <= SYNTHESIZED_WIRE_4(31);
ELSE
	gdfx_temp0(31) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(30) <= SYNTHESIZED_WIRE_4(30);
ELSE
	gdfx_temp0(30) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(29) <= SYNTHESIZED_WIRE_4(29);
ELSE
	gdfx_temp0(29) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(28) <= SYNTHESIZED_WIRE_4(28);
ELSE
	gdfx_temp0(28) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(27) <= SYNTHESIZED_WIRE_4(27);
ELSE
	gdfx_temp0(27) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(26) <= SYNTHESIZED_WIRE_4(26);
ELSE
	gdfx_temp0(26) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(25) <= SYNTHESIZED_WIRE_4(25);
ELSE
	gdfx_temp0(25) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(24) <= SYNTHESIZED_WIRE_4(24);
ELSE
	gdfx_temp0(24) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(23) <= SYNTHESIZED_WIRE_4(23);
ELSE
	gdfx_temp0(23) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(22) <= SYNTHESIZED_WIRE_4(22);
ELSE
	gdfx_temp0(22) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(21) <= SYNTHESIZED_WIRE_4(21);
ELSE
	gdfx_temp0(21) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(20) <= SYNTHESIZED_WIRE_4(20);
ELSE
	gdfx_temp0(20) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(19) <= SYNTHESIZED_WIRE_4(19);
ELSE
	gdfx_temp0(19) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(18) <= SYNTHESIZED_WIRE_4(18);
ELSE
	gdfx_temp0(18) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(17) <= SYNTHESIZED_WIRE_4(17);
ELSE
	gdfx_temp0(17) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(16) <= SYNTHESIZED_WIRE_4(16);
ELSE
	gdfx_temp0(16) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(15) <= SYNTHESIZED_WIRE_4(15);
ELSE
	gdfx_temp0(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(14) <= SYNTHESIZED_WIRE_4(14);
ELSE
	gdfx_temp0(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(13) <= SYNTHESIZED_WIRE_4(13);
ELSE
	gdfx_temp0(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(12) <= SYNTHESIZED_WIRE_4(12);
ELSE
	gdfx_temp0(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(11) <= SYNTHESIZED_WIRE_4(11);
ELSE
	gdfx_temp0(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(10) <= SYNTHESIZED_WIRE_4(10);
ELSE
	gdfx_temp0(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(9) <= SYNTHESIZED_WIRE_4(9);
ELSE
	gdfx_temp0(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(8) <= SYNTHESIZED_WIRE_4(8);
ELSE
	gdfx_temp0(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(7) <= SYNTHESIZED_WIRE_4(7);
ELSE
	gdfx_temp0(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(6) <= SYNTHESIZED_WIRE_4(6);
ELSE
	gdfx_temp0(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(5) <= SYNTHESIZED_WIRE_4(5);
ELSE
	gdfx_temp0(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(4) <= SYNTHESIZED_WIRE_4(4);
ELSE
	gdfx_temp0(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(3) <= SYNTHESIZED_WIRE_4(3);
ELSE
	gdfx_temp0(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(2) <= SYNTHESIZED_WIRE_4(2);
ELSE
	gdfx_temp0(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(1) <= SYNTHESIZED_WIRE_4(1);
ELSE
	gdfx_temp0(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_4,ALU_2_DBus_ALTERA_SYNTHESIZED)
BEGIN
if (ALU_2_DBus_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(0) <= SYNTHESIZED_WIRE_4(0);
ELSE
	gdfx_temp0(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(31) <= SYNTHESIZED_WIRE_5(31);
ELSE
	gdfx_temp0(31) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(30) <= SYNTHESIZED_WIRE_5(30);
ELSE
	gdfx_temp0(30) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(29) <= SYNTHESIZED_WIRE_5(29);
ELSE
	gdfx_temp0(29) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(28) <= SYNTHESIZED_WIRE_5(28);
ELSE
	gdfx_temp0(28) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(27) <= SYNTHESIZED_WIRE_5(27);
ELSE
	gdfx_temp0(27) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(26) <= SYNTHESIZED_WIRE_5(26);
ELSE
	gdfx_temp0(26) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(25) <= SYNTHESIZED_WIRE_5(25);
ELSE
	gdfx_temp0(25) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(24) <= SYNTHESIZED_WIRE_5(24);
ELSE
	gdfx_temp0(24) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(23) <= SYNTHESIZED_WIRE_5(23);
ELSE
	gdfx_temp0(23) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(22) <= SYNTHESIZED_WIRE_5(22);
ELSE
	gdfx_temp0(22) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(21) <= SYNTHESIZED_WIRE_5(21);
ELSE
	gdfx_temp0(21) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(20) <= SYNTHESIZED_WIRE_5(20);
ELSE
	gdfx_temp0(20) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(19) <= SYNTHESIZED_WIRE_5(19);
ELSE
	gdfx_temp0(19) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(18) <= SYNTHESIZED_WIRE_5(18);
ELSE
	gdfx_temp0(18) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(17) <= SYNTHESIZED_WIRE_5(17);
ELSE
	gdfx_temp0(17) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(16) <= SYNTHESIZED_WIRE_5(16);
ELSE
	gdfx_temp0(16) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(15) <= SYNTHESIZED_WIRE_5(15);
ELSE
	gdfx_temp0(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(14) <= SYNTHESIZED_WIRE_5(14);
ELSE
	gdfx_temp0(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(13) <= SYNTHESIZED_WIRE_5(13);
ELSE
	gdfx_temp0(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(12) <= SYNTHESIZED_WIRE_5(12);
ELSE
	gdfx_temp0(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(11) <= SYNTHESIZED_WIRE_5(11);
ELSE
	gdfx_temp0(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(10) <= SYNTHESIZED_WIRE_5(10);
ELSE
	gdfx_temp0(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(9) <= SYNTHESIZED_WIRE_5(9);
ELSE
	gdfx_temp0(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(8) <= SYNTHESIZED_WIRE_5(8);
ELSE
	gdfx_temp0(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(7) <= SYNTHESIZED_WIRE_5(7);
ELSE
	gdfx_temp0(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(6) <= SYNTHESIZED_WIRE_5(6);
ELSE
	gdfx_temp0(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(5) <= SYNTHESIZED_WIRE_5(5);
ELSE
	gdfx_temp0(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(4) <= SYNTHESIZED_WIRE_5(4);
ELSE
	gdfx_temp0(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(3) <= SYNTHESIZED_WIRE_5(3);
ELSE
	gdfx_temp0(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(2) <= SYNTHESIZED_WIRE_5(2);
ELSE
	gdfx_temp0(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(1) <= SYNTHESIZED_WIRE_5(1);
ELSE
	gdfx_temp0(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(SYNTHESIZED_WIRE_5,SYNTHESIZED_WIRE_6)
BEGIN
if (SYNTHESIZED_WIRE_6 = '1') THEN
	gdfx_temp0(0) <= SYNTHESIZED_WIRE_5(0);
ELSE
	gdfx_temp0(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(31) <= IO_IN(31);
ELSE
	gdfx_temp0(31) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(30) <= IO_IN(30);
ELSE
	gdfx_temp0(30) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(29) <= IO_IN(29);
ELSE
	gdfx_temp0(29) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(28) <= IO_IN(28);
ELSE
	gdfx_temp0(28) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(27) <= IO_IN(27);
ELSE
	gdfx_temp0(27) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(26) <= IO_IN(26);
ELSE
	gdfx_temp0(26) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(25) <= IO_IN(25);
ELSE
	gdfx_temp0(25) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(24) <= IO_IN(24);
ELSE
	gdfx_temp0(24) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(23) <= IO_IN(23);
ELSE
	gdfx_temp0(23) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(22) <= IO_IN(22);
ELSE
	gdfx_temp0(22) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(21) <= IO_IN(21);
ELSE
	gdfx_temp0(21) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(20) <= IO_IN(20);
ELSE
	gdfx_temp0(20) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(19) <= IO_IN(19);
ELSE
	gdfx_temp0(19) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(18) <= IO_IN(18);
ELSE
	gdfx_temp0(18) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(17) <= IO_IN(17);
ELSE
	gdfx_temp0(17) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(16) <= IO_IN(16);
ELSE
	gdfx_temp0(16) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(15) <= IO_IN(15);
ELSE
	gdfx_temp0(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(14) <= IO_IN(14);
ELSE
	gdfx_temp0(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(13) <= IO_IN(13);
ELSE
	gdfx_temp0(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(12) <= IO_IN(12);
ELSE
	gdfx_temp0(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(11) <= IO_IN(11);
ELSE
	gdfx_temp0(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(10) <= IO_IN(10);
ELSE
	gdfx_temp0(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(9) <= IO_IN(9);
ELSE
	gdfx_temp0(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(8) <= IO_IN(8);
ELSE
	gdfx_temp0(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(7) <= IO_IN(7);
ELSE
	gdfx_temp0(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(6) <= IO_IN(6);
ELSE
	gdfx_temp0(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(5) <= IO_IN(5);
ELSE
	gdfx_temp0(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(4) <= IO_IN(4);
ELSE
	gdfx_temp0(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(3) <= IO_IN(3);
ELSE
	gdfx_temp0(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(2) <= IO_IN(2);
ELSE
	gdfx_temp0(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(1) <= IO_IN(1);
ELSE
	gdfx_temp0(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(IO_IN,IO_2_Reg_ALTERA_SYNTHESIZED)
BEGIN
if (IO_2_Reg_ALTERA_SYNTHESIZED = '1') THEN
	gdfx_temp0(0) <= IO_IN(0);
ELSE
	gdfx_temp0(0) <= 'Z';
END IF;
END PROCESS;


PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(31) <= Rs1(31);
ELSE
	IO_OUT(31) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(30) <= Rs1(30);
ELSE
	IO_OUT(30) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(29) <= Rs1(29);
ELSE
	IO_OUT(29) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(28) <= Rs1(28);
ELSE
	IO_OUT(28) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(27) <= Rs1(27);
ELSE
	IO_OUT(27) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(26) <= Rs1(26);
ELSE
	IO_OUT(26) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(25) <= Rs1(25);
ELSE
	IO_OUT(25) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(24) <= Rs1(24);
ELSE
	IO_OUT(24) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(23) <= Rs1(23);
ELSE
	IO_OUT(23) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(22) <= Rs1(22);
ELSE
	IO_OUT(22) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(21) <= Rs1(21);
ELSE
	IO_OUT(21) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(20) <= Rs1(20);
ELSE
	IO_OUT(20) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(19) <= Rs1(19);
ELSE
	IO_OUT(19) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(18) <= Rs1(18);
ELSE
	IO_OUT(18) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(17) <= Rs1(17);
ELSE
	IO_OUT(17) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(16) <= Rs1(16);
ELSE
	IO_OUT(16) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(15) <= Rs1(15);
ELSE
	IO_OUT(15) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(14) <= Rs1(14);
ELSE
	IO_OUT(14) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(13) <= Rs1(13);
ELSE
	IO_OUT(13) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(12) <= Rs1(12);
ELSE
	IO_OUT(12) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(11) <= Rs1(11);
ELSE
	IO_OUT(11) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(10) <= Rs1(10);
ELSE
	IO_OUT(10) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(9) <= Rs1(9);
ELSE
	IO_OUT(9) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(8) <= Rs1(8);
ELSE
	IO_OUT(8) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(7) <= Rs1(7);
ELSE
	IO_OUT(7) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(6) <= Rs1(6);
ELSE
	IO_OUT(6) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(5) <= Rs1(5);
ELSE
	IO_OUT(5) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(4) <= Rs1(4);
ELSE
	IO_OUT(4) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(3) <= Rs1(3);
ELSE
	IO_OUT(3) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(2) <= Rs1(2);
ELSE
	IO_OUT(2) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(1) <= Rs1(1);
ELSE
	IO_OUT(1) <= 'Z';
END IF;
END PROCESS;

PROCESS(Rs1,Reg_2_IO_ALTERA_SYNTHESIZED)
BEGIN
if (Reg_2_IO_ALTERA_SYNTHESIZED = '1') THEN
	IO_OUT(0) <= Rs1(0);
ELSE
	IO_OUT(0) <= 'Z';
END IF;
END PROCESS;


b2v_UC : uc
PORT MAP(clear => reset,
		 clock => clock,
		 instruction => instruction_ALTERA_SYNTHESIZED(31 DOWNTO 29),
		 IR_Ld => IR_Ld_ALTERA_SYNTHESIZED,
		 PC_Inc => Pc_Inc_ALTERA_SYNTHESIZED,
		 ALU_2_DBus => ALU_2_DBus_ALTERA_SYNTHESIZED,
		 DM_Rd => DM_Rd_ALTERA_SYNTHESIZED,
		 DM_Wr => DM_Wr_ALTERA_SYNTHESIZED,
		 PC_Ld_En => PC_Ld_En_ALTERA_SYNTHESIZED,
		 Reg_2_IO => Reg_2_IO_ALTERA_SYNTHESIZED,
		 IO_2_Reg => IO_2_Reg_ALTERA_SYNTHESIZED,
		 Reg_Wr => Reg_Wr_ALTERA_SYNTHESIZED,
		 Stat_Wr => Stat_Wr_ALTERA_SYNTHESIZED,
		 DM_2_DBus => DM_2_DBus_ALTERA_SYNTHESIZED);

Pc_Ld <= Pc_Ld_ALTERA_SYNTHESIZED;
IR_Ld <= IR_Ld_ALTERA_SYNTHESIZED;
Pc_Inc <= Pc_Inc_ALTERA_SYNTHESIZED;
ALU_2_DBus <= ALU_2_DBus_ALTERA_SYNTHESIZED;
DM_Rd <= DM_Rd_ALTERA_SYNTHESIZED;
DM_Wr <= DM_Wr_ALTERA_SYNTHESIZED;
PC_Ld_En <= PC_Ld_En_ALTERA_SYNTHESIZED;
Reg_2_IO <= Reg_2_IO_ALTERA_SYNTHESIZED;
IO_2_Reg <= IO_2_Reg_ALTERA_SYNTHESIZED;
Reg_Wr <= Reg_Wr_ALTERA_SYNTHESIZED;
Stat_Wr <= Stat_Wr_ALTERA_SYNTHESIZED;
DM_2_DBus <= DM_2_DBus_ALTERA_SYNTHESIZED;
DBus <= gdfx_temp0;
IM_address <= addr;
IM_instruction_out <= preir;
instruction <= instruction_ALTERA_SYNTHESIZED;
RSource1 <= Rs1;
RSource2 <= Rs2;
stat_CVNZ(3 DOWNTO 0) <= stat(3 DOWNTO 0);

gnd <= '0';
vcc <= '1';
END bdf_type;